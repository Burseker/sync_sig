--=============================
-- Developed by SVB. Ver. 0.2.0 
--=============================
----------------------------------------------------------------------------------
-- Company:         ������-�����
-- Engineer:        ������ �������
--                  
-- Create Date:     18.03.2014
-- Design Name:     pckr8to32
-- Module Name:     pckr8to32 - Beh
-- Project Name:    Quartet
-- Target Devices:  Stratix II: EP2S60F484I4
-- Tool versions:   Notepad++
-- Description:     ����������� ��������� ������ �� 8� � 32�
--                  �������� ���
--                  
--                  
-- Dependencies:    
--                  
-- Revision:        
-- Revision 0.0.0 - File created   
-- Revision 0.1.0 - ��������� ���� �� pckr8to16 � pckr16to18
-- Revision 0.2.0 - �������� �������� ����������� ENDIANNESS
--
--                  
-- Additional Comments: 
-- 
--     
-- 
-- 
-- 
-- 
-- 
----------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use work.pkg_sim.all;
use work.pkg_func.all;
--=========================

entity pckr8to32 is
    generic(
        ENDIANNESS : string := "BIG_ENDIAN" -- "BIG_ENDIAN", "LITTLE_ENDIAN"
    );
    port (
        aclr    : in  std_logic;
        clk     : in  std_logic;
        
        idat    : in  std_logic_vector(7 downto 0);
        istb    : in  std_logic;
        iend    : in  std_logic;
        iten    : out std_logic;
        
        odat    : out std_logic_vector(31 downto 0);
        ostb    : out std_logic;
        oend    : out std_logic;
        oten    : in  std_logic
    );
end pckr8to32;

architecture beh of pckr8to32 is

    constant C_IWIDTH   : natural := 8;
    constant C_OWIDTH   : natural := 32;
    
    signal s_iten        : std_logic := '0';
    
    signal s_adat        : std_logic_vector( 15 downto 0) := (others => '0');
    signal s_aend        : std_logic := '0';
    signal s_astb        : std_logic := '0';
    signal s_aten        : std_logic := '0';
    
    signal s_odat        : std_logic_vector( C_OWIDTH-1 downto 0) := (others => '0');
    signal s_oend        : std_logic := '0';
    signal s_ostb        : std_logic := '0';
    
begin
    
--=============================================
-- TYPICAL PROCESS
--=============================================
    -- process(aclr, clk)
    -- begin
        -- if(aclr = '1')then
        -- elsif(rising_edge(clk))then
        -- end if;
    -- end process;
    
    
--=============================================
--���������� ������� � 16
--=============================================
pckr8to16inst: entity work.pckr8to16
generic map( ENDIANNESS => ENDIANNESS)
port map(
    aclr    => aclr,
    clk     => clk,
    
    idat    => idat,
    istb    => istb,
    iend    => iend,
    iten    => s_iten,
    
    odat    => s_adat,
    ostb    => s_astb,
    oend    => s_aend,
    oten    => s_aten
);


--=============================================
--���������� ������� � 18
--=============================================
pckr16to18inst: entity work.pckr16to32
generic map( ENDIANNESS => ENDIANNESS)
port map(
    aclr    => aclr,
    clk     => clk,
    
    idat    => s_adat,
    istb    => s_astb,
    iend    => s_aend,
    iten    => s_aten,
    
    odat    => s_odat,
    ostb    => s_ostb,
    oend    => s_oend,
    oten    => oten
);


--==================================
-- ���������� �������� ��������
--==================================   
    iten <= s_iten;
    
    odat <= s_odat;
    ostb <= s_ostb;
    oend <= s_oend;
    
end Beh;
